module main;
initial begin
	$display("main");
	$finish;
end
endmodule

module top;
initial begin
	$display("top");
	$finish;
end
endmodule
